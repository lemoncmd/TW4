module cpu (
    input logic clock,
    input logic reset,
    output logic [5:0] addr,
    input logic [7:0] data,
    input logic [3:0] in,
    output logic [3:0] out
);

endmodule

